library verilog;
use verilog.vl_types.all;
entity img_processing_tb is
end img_processing_tb;
