library verilog;
use verilog.vl_types.all;
entity number_display_vlg_vec_tst is
end number_display_vlg_vec_tst;
